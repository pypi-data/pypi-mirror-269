Begin3
Language:    SV, 850
Title:       GNU chcp-typsnitt
Description: LOADFONT (GNUCHCP) r�a EGA-/VGA-bitmappstypsnitt f�r textl�gen.
Keywords:    loadfont gnuchcp bitmapp typsnitt ega vga sk�rm
End
